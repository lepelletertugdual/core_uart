-- #################################################################################################################################################################################
-- file :
--     core_uart_tx.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     UART receiver
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     register tranfer level (RTL)
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     clock ratio must be higher or equal to 16.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2024-04-25
--         file creation
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--     02. entity
--     03. architecture
--         03.01. constants
--         03.02. signals
--         03.03. input assignment
--         03.04. alive output pin generation
--         03.05. output assignment
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;

    -- =============================================================================================================================================================================
	-- 01.01. custom
    -- =============================================================================================================================================================================	
	library work;
	    use work.pkg_core_uart_rx.all;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity core_uart_rx is
    generic (
	     g_clk_i_freq  : integer := 100_000_000
		;g_baud        : integer :=     115_200
		;g_data_length : integer :=           8
	);
    port (
	     i_clk     : in  std_logic
		;i_rst     : in  std_logic
		;o_data_en : out std_logic
		;o_data    : out std_logic_vector(g_data_length-1 downto 0)
		;o_ready   : out std_logic
		;o_done    : out std_logic
		;i_rx      : in  std_logic
		;o_error   : out std_logic_vector(7 downto 0)
	);
end entity core_uart_rx;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture rtl of core_uart_rx is

    -- =============================================================================================================================================================================
	-- 03.01. constants
    -- =============================================================================================================================================================================
	constant c_over_sampling : integer := 16;
    constant c_clk_ratio     : integer := integer(real(g_clk_i_freq)/(real(c_over_sampling)*real(g_baud)));

    -- =============================================================================================================================================================================
	-- 03.04. types
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. FSM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        type t_fsm_main is (
		     state_fsm_main_idle
		    ,state_fsm_main_start
			,state_fsm_main_data
			,state_fsm_main_stop
		);
	
    -- =============================================================================================================================================================================
	-- 03.02. signals
    -- =============================================================================================================================================================================
	signal s_clk           : std_logic;
	signal s_rst           : std_logic;
	signal s_error_ratio   : std_logic;
	signal s_data          : std_logic_vector(g_data_length-1 downto 0);
	signal s_data_en       : std_logic;
	signal s_data_reg      : std_logic_vector(g_data_length-1 downto 0);
	signal s_cnt_bit       : integer range 0 to g_data_length-1;
	signal s_rx            : std_logic;
	signal s_ready         : std_logic;
	signal s_done          : std_logic;
	signal s_tick          : std_logic;
	signal s_rx_meta       : std_logic;
	signal s_rx_sync       : std_logic;
	signal s_cnt_baud_rate : integer range 0 to c_clk_ratio-1;
	signal s_cnt_tick      : integer range 0 to c_over_sampling-1;
	signal s_fsm_main      : t_fsm_main;
	
begin
    -- =============================================================================================================================================================================
	-- 03.03. check input parameters
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. check clock ratio
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    check_clk_ratio_ok : if (c_clk_ratio > c_clk_ratio_upper_bound or c_clk_ratio = c_clk_ratio_upper_bound) generate
	        s_error_ratio <= '0';
	    end generate check_clk_ratio_ok;

	    check_clk_ratio_ko : if (c_clk_ratio < c_clk_ratio_upper_bound) generate
	        s_error_ratio <= '1';
	    end generate check_clk_ratio_ko;

    -- =============================================================================================================================================================================
	-- 03.04. input assignment
    -- =============================================================================================================================================================================
	s_clk     <= i_clk;
	s_rst     <= i_rst;
    s_rx      <= i_rx;

    -- =============================================================================================================================================================================
	-- 03.05. baud rate generator
    -- =============================================================================================================================================================================
    p_gen_baud_rate : process(s_clk,s_rst)
	begin
	    if (s_rst = '1') then
		    s_cnt_baud_rate <= 0;
			s_tick <= '0';
		elsif (rising_edge(s_clk)) then
		    s_tick <= '0';
		    if (s_cnt_baud_rate = c_clk_ratio-1) then
			    s_cnt_baud_rate <= 0;
				s_tick <= '1';
            else
			    s_cnt_baud_rate <= s_cnt_baud_rate + 1;
			end if;
		end if;
	end process p_gen_baud_rate;

    -- =============================================================================================================================================================================
	-- 03.05. resynchronization stage
    -- =============================================================================================================================================================================
    p_resync_rx : process(s_clk,s_rst)
	begin
	    if (s_rst = '1') then
		    s_rx_meta <= '1';
			s_rx_sync <= '1';
		elsif (rising_edge(s_clk)) then
		    s_rx_meta <= s_rx;
			s_rx_sync <= s_rx_meta;
		end if;
	end process p_resync_rx;

    -- =============================================================================================================================================================================
	-- 03.05. main FSM
    -- =============================================================================================================================================================================
    p_fsm_main : process(s_clk,s_rst)
	begin
	    if (s_rst = '1') then
		    s_ready <= '0';
			s_done <= '0';
			s_data_en <= '0';
			s_data <= (others => '0');
		    s_data_reg <= (others => '0');
			s_fsm_main <= state_fsm_main_idle;
		elsif (rising_edge(s_clk)) then
		    s_done <= '0';
		    case s_fsm_main is
			    when state_fsm_main_idle =>
				    s_ready <= '1';
				    -- detection start bit
				    if (s_rx_sync = '0') then
					    s_ready <= '0';
						s_data_en <= '0';
					    s_fsm_main <= state_fsm_main_start;
					end if;
				when state_fsm_main_start =>
				    -- detection baud rate tick
				    if (s_tick = '1') then
					    -- reach middle start bit
					    if (s_cnt_tick = c_over_sampling/2-1) then
						    s_cnt_tick <= 0;
							s_fsm_main <= state_fsm_main_data;
						else
						    s_cnt_tick <= s_cnt_tick + 1;
						end if;
					end if;
				when state_fsm_main_data  =>
				    -- detection baud rate tick
				    if (s_tick = '1') then
					    -- reach middle data bit
					    if (s_cnt_tick = c_over_sampling-1) then
						    s_cnt_tick <= 0;
							-- sample rx data bit
							s_data_reg <= s_data_reg(s_data_reg'length-2 downto 0) & s_rx_sync;
							-- process all data bits
							if (s_cnt_bit = g_data_length-1) then
							    s_cnt_bit <= 0;
							    s_fsm_main <= state_fsm_main_stop;
                            else
							    s_cnt_bit <= s_cnt_bit + 1;
							end if;
						else
						    s_cnt_tick <= s_cnt_tick + 1;
						end if;
					else
					end if;
				when state_fsm_main_stop  =>
				    -- detection baud rate tick
				    if (s_tick = '1') then
					    -- reach middle start bit
					    if (s_cnt_tick = c_over_sampling-1) then
						    s_cnt_tick <= 0;
							s_ready <= '1';
							s_done <= '1';
							s_data_en <= '1';
							s_data <= s_data_reg;
							s_fsm_main <= state_fsm_main_idle;
						else
						    s_cnt_tick <= s_cnt_tick + 1;
						end if;
					end if;
			end case;
		end if;
	end process p_fsm_main;

    -- =============================================================================================================================================================================
	-- 03.06. output assignment
    -- =============================================================================================================================================================================
	o_done    <= s_done;
	o_ready   <= s_ready;
	o_data    <= s_data;
	o_data_en <= s_data_en;
    o_error   <= (
	     c_pos_error_ratio => s_error_ratio
		,others            => '0'
	);

end architecture rtl;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################