-- #################################################################################################################################################################################
-- file :
--     core_uart_tx.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     UART transmitter
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     register tranfer level (RTL)
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     clock ratio must be higher or equal to 16.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2024-04-23
--         file creation
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--     02. entity
--     03. architecture
--         03.01. constants
--         03.02. signals
--         03.03. input assignment
--         03.04. alive output pin generation
--         03.05. output assignment
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity core_uart is
    generic (
	     g_clk_i_freq  : integer := 100_000_000
		;g_baud        : integer :=     115_200
		;g_data_length : integer :=           8
	);
    port (
	     i_clk        : in  std_logic
		;i_rst        : in  std_logic
		-- transmitter
		;i_tx_data_en : in  std_logic
		;i_tx_data    : in  std_logic_vector(g_data_length-1 downto 0)
		;o_tx_ready   : out std_logic
		;o_tx_done    : out std_logic
		;o_tx_line    : out std_logic
		;o_tx_error   : out std_logic_vector(7 downto 0)
		-- receiver
		;o_rx_data_en : out std_logic
		;o_rx_data    : out std_logic_vector(g_data_length-1 downto 0)
		;o_rx_ready   : out std_logic
		;o_rx_done    : out std_logic
		;i_rx_line    : in  std_logic
		;o_rx_error   : out std_logic_vector(7 downto 0)
	);
end entity core_uart;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture schematic of core_uart is

    -- =============================================================================================================================================================================
	-- 03.01. component declaration
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. core_uart_rx
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component core_uart_rx is
            generic (
	             g_clk_i_freq  : integer := 100_000_000
		        ;g_baud        : integer :=     115_200
		        ;g_data_length : integer :=           8
	        );
            port (
	             i_clk     : in  std_logic
		        ;i_rst     : in  std_logic
		        ;o_data_en : out std_logic
		        ;o_data    : out std_logic_vector(g_data_length-1 downto 0)
		        ;o_ready   : out std_logic
		        ;o_done    : out std_logic
		        ;i_rx      : in  std_logic
		        ;o_error   : out std_logic_vector(7 downto 0)
	        );
        end component core_uart_rx;
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. core_uart_rx
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    component core_uart_tx is
            generic (
	             g_clk_i_freq  : integer := 100_000_000
		        ;g_baud        : integer :=     115_200
		        ;g_data_length : integer :=           8
	        );
            port (
	             i_clk     : in  std_logic
		        ;i_rst     : in  std_logic
		        ;i_data_en : in  std_logic
		        ;i_data    : in  std_logic_vector(g_data_length-1 downto 0)
		        ;o_ready   : out std_logic
		        ;o_done    : out std_logic
		        ;o_tx      : out std_logic
		        ;o_error   : out std_logic_vector(7 downto 0)
	        );
        end component core_uart_tx;
	
    -- =============================================================================================================================================================================
	-- 03.01. signal declaration
    -- =============================================================================================================================================================================
    signal s_clk        : std_logic;
	signal s_rst        : std_logic;
	signal s_tx_data_en : std_logic;
	signal s_tx_data    : std_logic_vector(g_data_length-1 downto 0);
	signal s_tx_ready   : std_logic;
	signal s_tx_done    : std_logic;
	signal s_tx_line    : std_logic;
	signal s_tx_error   : std_logic_vector(7 downto 0);
	signal s_rx_data_en : std_logic;
	signal s_rx_data    : std_logic_vector(g_data_length-1 downto 0);
	signal s_rx_ready   : std_logic;
	signal s_rx_done    : std_logic;
	signal s_rx_line    : std_logic;
	signal s_rx_error   : std_logic_vector(7 downto 0);
	
begin
 
    -- =============================================================================================================================================================================
	-- 03.04. input assignment
    -- =============================================================================================================================================================================
    s_clk <= i_clk;            
	s_rst <= i_rst;
	s_tx_data_en <= i_tx_data_en;
	s_tx_data <= i_tx_data;     
	s_rx_line <= i_rx_line;    

    -- =============================================================================================================================================================================
	-- 03.04. component instanciation
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. core_uart_tx
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    inst_core_uart_tx : core_uart_tx
            generic map (
	             g_clk_i_freq  => g_clk_i_freq
	            ,g_baud        => g_baud
	            ,g_data_length => g_data_length
	        )
            port map (
	             i_clk     => s_clk
	            ,i_rst     => s_rst
	            ,i_data_en => s_tx_data_en 
	            ,i_data    => s_tx_data
	            ,o_ready   => s_tx_ready
	            ,o_done    => s_tx_done
	            ,o_tx      => s_tx_line
	            ,o_error   => s_tx_error
	        );

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. core_uart_rx
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_core_uart_rx : core_uart_rx
            generic map (
	             g_clk_i_freq  => g_clk_i_freq
		        ,g_baud        => g_baud
		        ,g_data_length => g_data_length
	        )
            port map (
	             i_clk     => s_clk
		        ,i_rst     => s_rst
		        ,o_data_en => s_rx_data_en
		        ,o_data    => s_rx_data
		        ,o_ready   => s_rx_ready
		        ,o_done    => s_rx_done
		        ,i_rx      => s_rx_line
		        ,o_error   => s_rx_error
	        );

    -- =============================================================================================================================================================================
	-- 03.04. output assignment
    -- =============================================================================================================================================================================
	o_tx_ready   <= s_tx_ready;
	o_tx_done    <= s_tx_done;
	o_tx_line    <= s_tx_line;
	o_tx_error   <= s_tx_error;
	o_rx_data_en <= s_rx_data_en;
	o_rx_data    <= s_rx_data;
	o_rx_ready   <= s_rx_ready;
	o_rx_done    <= s_rx_done;
	o_rx_error   <= s_rx_error;
	
end architecture schematic;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################