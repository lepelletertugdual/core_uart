-- #################################################################################################################################################################################
-- file :
--     bch_core_uart.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     core_uart.vhd testbench file.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     behavioral
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     none
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2023-11-11
--         file creation
--     2024-10-28
--         changing the host clock frequency and adaptating the testbench to manage three clock domains
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
-- 01. libraries
--    01.01. standard
--	  01.02. custom
-- 02. entity
-- 03. architecture
    -- 03.01. component declaration
	    -- 03.01.01. DUT : core_uart
	-- 03.02. files
	    -- 03.02.01. LOG
		-- 03.02.02. RPT
	-- 03.03. types
	    -- 03.03.01. FSM
		    -- 03.03.01.01. fsm_main
			-- 03.03.01.02. fsm_init
			-- 03.03.01.03. fsm_test
			-- 03.03.01.04. fsm_file_mgt_log
			-- 03.03.01.05. fsm_file_mgt_rpt
		-- 03.03.02. test status
		-- 03.03.03. array
	-- 03.04. constants
	    -- 03.04.01. SIM
		-- 03.04.02. oscillator
		-- 03.04.03. DUT : core_uart
		-- 03.04.04. HOST
		-- 03.04.05. clocks ratios
		-- 03.04.06. files
	-- 03.05. signals
	    -- 03.05.01. SIM
		    -- 03.05.01.01. FSM
			-- 03.05.01.02. files
			-- 03.05.01.03. clocks
			-- 03.05.01.04. reset
			-- 03.05.01.05. testbench
		-- 03.05.02. DUT : core_uart
		    -- 03.05.02.01. clock
			-- 03.05.02.02. reset
			-- 03.05.02.03. core_uart_tx
			-- 03.05.02.04. core_uart_rx
		-- 03.05.03. HOST
		    -- 03.05.03.01. clock
			-- 03.05.03.02. reset
			-- 03.05.03.03. core_uart_tx
			-- 03.05.03.04. core_uart_rx
	-- 03.06. reset management
	    -- 03.06.01. SIM
		-- 03.06.02. DUT
		-- 03.06.03. HOST
	-- 03.07. clock generation
	    -- 03.07.01. SIM
		-- 03.07.02. oscillator
		-- 03.07.03. HOST
	-- 03.08. clock assignment
	-- 03.09. component instantiation
	    -- 03.09.01. HOST : core_uart
		-- 03.09.02. loopback
		-- 03.09.03. DUT : core_uart
	-- 03.10. clock domain crossing (CDC)
	    -- 03.10.01. from SIM to DUT (from fast to slow)
		-- 03.10.02. from SIM to HST (from fast to slow)
		-- 03.10.03. edge detector from HST to SIM (from slow to fast)
		-- 03.10.04. edge detector from DUT to SIM (from slow to fast)
	-- 03.11. fsm_main
	-- 03.12. fsm_init
	-- 03.13. fsm_test
	-- 03.14. fsm_file_mgt_log
	-- 03.15. fsm_file_mgt_rpt
	-- 03.16. error detection
	-- 03.17. simulation abort
	-- 03.18. end of simulation
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;
	
    library std;
        use std.textio.all;

    -- =============================================================================================================================================================================
	-- 01.02. custom
    -- =============================================================================================================================================================================
    library work;
        use work.pkg_mgt_file.all;
		use work.pkg_core_uart_tx.all;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity bch_core_uart is
end entity bch_core_uart;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture behavioral of bch_core_uart is

    -- =============================================================================================================================================================================
	-- 03.01. component declaration
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. DUT : core_uart
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component core_uart is
            generic (
	         g_clk_i_freq  : integer := 100_000_000
		    ;g_baud        : integer :=     115_200
		    ;g_data_length : integer :=           8
	    );
        port (
	         i_clk        : in  std_logic
		    ;i_rst        : in  std_logic
		    -- transmitter
		    ;i_tx_data_en : in  std_logic
		    ;i_tx_data    : in  std_logic_vector(g_data_length-1 downto 0)
		    ;o_tx_ready   : out std_logic
		    ;o_tx_done    : out std_logic
		    ;o_tx_line    : out std_logic
		    ;o_tx_error   : out std_logic_vector(7 downto 0)
		    -- receiver
		    ;o_rx_data_en : out std_logic
		    ;o_rx_data    : out std_logic_vector(g_data_length-1 downto 0)
		    ;o_rx_ready   : out std_logic
		    ;o_rx_done    : out std_logic
		    ;i_rx_line    : in  std_logic
		    ;o_rx_error   : out std_logic_vector(7 downto 0)
	    );
        end component core_uart;

    -- =============================================================================================================================================================================
	-- 03.02. files
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.01. LOG
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_log : text;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.02. RPT
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_rpt : text;

    -- =============================================================================================================================================================================
	-- 03.03. types
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. FSM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.03.01.01. fsm_main
			-- =====================================================================================================================================================================
	        type t_fsm_main is (
	             state_fsm_main_start
                ,state_fsm_main_file_rpt_open
                ,state_fsm_main_file_log_open
			    ,state_fsm_main_init
		        ,state_fsm_main_run
                ,state_fsm_main_file_rpt_close
                ,state_fsm_main_file_log_close
		        ,state_fsm_main_stop
	        );

		    -- =====================================================================================================================================================================
			-- 03.03.01.02. fsm_init
			-- =====================================================================================================================================================================
	        type t_fsm_init is (
	             state_fsm_init_idle
		        ,state_fsm_init_run
		        ,state_fsm_init_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.03.01.03. fsm_test
			-- =====================================================================================================================================================================
	        type t_fsm_test is (
	             state_fsm_test_idle
				,state_fsm_test_dut_to_hst_send_data
		        ,state_fsm_test_dut_to_hst_wait_ready
		        ,state_fsm_test_dut_to_hst_wait_done
				,state_fsm_test_dut_to_hst_check_data
				,state_fsm_test_hst_to_dut_send_data
		        ,state_fsm_test_hst_to_dut_wait_ready
		        ,state_fsm_test_hst_to_dut_wait_done
				,state_fsm_test_hst_to_dut_check_data
				,state_fsm_test_done
	        );
	
		    -- =====================================================================================================================================================================
			-- 03.03.01.04. fsm_file_mgt_log
			-- =====================================================================================================================================================================
	        type t_fsm_file_mgt_log is (
	             state_fsm_file_mgt_log_open
				,state_fsm_file_mgt_log_write_head
	            ,state_fsm_file_mgt_log_write_data
		        ,state_fsm_file_mgt_log_close
				,state_fsm_file_mgt_log_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.03.01.05. fsm_file_mgt_rpt
			-- =====================================================================================================================================================================
	        type t_fsm_file_mgt_rpt is (
	             state_fsm_file_mgt_rpt_open
	            ,state_fsm_file_mgt_rpt_write_status
		        ,state_fsm_file_mgt_rpt_close
				,state_fsm_file_mgt_rpt_done
	        );

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.02. test status
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	        type t_sim_test_status is (
	             TEST_OK
	            ,TEST_KO
	        );
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.03. array
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        type t_array_data is array (natural range <>) of std_logic_vector(7 downto 0);

    -- =============================================================================================================================================================================
	-- 03.04. constants
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_sim_clk_freq      : integer := 1_000_000_000;
	    constant c_sim_clk_delay     : time    := 0.9 us;
	    constant c_sim_rst_delay     : time    := 0.3 us;
        constant c_sim_clk_period_ns : time    := integer((real(1)/real(c_sim_clk_freq))*1.0e9)*1 ns;
	    constant c_sim_clk_period    : real    := real(1)/real(c_sim_clk_freq);	

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.02. oscillator
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_osc_delay     : time := 2.4 us;
	    constant c_osc_freq      : integer := 100_000_000;
        constant c_osc_period_ns : time := integer((real(1)/real(c_osc_freq))*1.0e9)*1 ns;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.03. DUT : core_uart
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_dut_rst_delay     : time    := 2.5 us;
	    constant c_dut_clk_freq      : integer := c_osc_freq;
		constant c_dut_clk_period    : real    := real(1)/real(c_dut_clk_freq);
		constant c_dut_baud          : integer := 115200;
		constant c_dut_data_length   : integer := 8;
	    constant c_array_data_length : integer := 2;
		constant c_array_data        : t_array_data(0 to c_array_data_length-1) := (
			    0 => x"A5",
				1 => x"5A"
			);
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.04. HOST
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        constant c_hst_clk_freq      : integer := 500_000_000;
		constant c_hst_clk_delay     : time    := 1.7 us;
	    constant c_hst_rst_delay     : time    := 5.7 us;
        constant c_hst_clk_period_ns : time    := integer((real(1)/real(c_hst_clk_freq))*1.0e9)*1 ns;
		constant c_hst_clk_period    : real    := real(1)/real(c_hst_clk_freq);
		constant c_hst_baud          : integer := 115200;
		constant c_hst_data_length   : integer := 8;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.05. clock ratios
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_ratio_clk_sim_clk_dut : integer := integer(real(c_sim_clk_freq)/real(c_dut_clk_freq));
		constant c_ratio_clk_sim_clk_hst : integer := integer(real(c_sim_clk_freq)/real(c_hst_clk_freq));
		
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.06. files
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_file_log_name : string := "log_bch_core_uart_wrapper_zedboard_sim.csv";
		constant c_file_rpt_name : string := "rpt_bch_core_uart_wrapper_zedboard_sim.txt";
	
    -- =============================================================================================================================================================================
	-- 03.05. signals
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.05.01.01. FSM
			-- =====================================================================================================================================================================
	        signal s_fsm_main_state   : t_fsm_main;
	        signal s_fsm_init_state   : t_fsm_init;
	        signal s_fsm_test_state   : t_fsm_test;
		    signal s_fsm_file_mgt_log : t_fsm_file_mgt_log;
		    signal s_fsm_file_mgt_rpt : t_fsm_file_mgt_rpt;
	
		    -- =====================================================================================================================================================================
			-- 03.05.01.02. files
			-- =====================================================================================================================================================================
		    signal s_sim_file_req_log_open  : std_logic;
		    signal s_sim_file_ack_log_open  : std_logic;
		    signal s_sim_file_req_log_close : std_logic;
		    signal s_sim_file_ack_log_close : std_logic;
		    signal s_sim_file_req_rpt_open  : std_logic;
		    signal s_sim_file_ack_rpt_open  : std_logic;
		    signal s_sim_file_req_rpt_close : std_logic;
		    signal s_sim_file_ack_rpt_close : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.01.03. clocks
			-- =====================================================================================================================================================================
            signal s_sim_clk : std_logic;
	        signal s_osc     : std_logic;
			signal s_hst_clk : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.01.04. reset
			-- =====================================================================================================================================================================
		    signal s_sim_rst : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.01.05. testbench
			-- =====================================================================================================================================================================
		    signal s_sim_done        : std_logic;
		    signal s_sim_init_req    : std_logic;
		    signal s_sim_init_ack    : std_logic;
		    signal s_sim_test_req    : std_logic;
		    signal s_sim_test_ack    : std_logic;
		    signal s_sim_test_status : t_sim_test_status;
			signal s_error           : std_logic;
			signal s_array_data_cnt  : integer range 0 to 1;
	        signal s_error_test      : std_logic;
			
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.02. DUT : core_uart
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.05.02.01. clock
			-- =====================================================================================================================================================================
            signal s_dut_i_clk : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.02. reset
			-- =====================================================================================================================================================================
	        signal s_dut_i_rst : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.03. core_uart_tx
			-- =====================================================================================================================================================================			
		    signal s_dut_uart_tx_i_data_en             : std_logic;
		    signal s_dut_uart_tx_i_data_en_reg         : std_logic_vector(c_ratio_clk_sim_clk_dut-1 downto 0);
			signal s_dut_uart_tx_i_data_en_reg_gen_tmp : std_logic_vector(c_ratio_clk_sim_clk_dut-1 downto 0);
			signal s_dut_uart_tx_i_data_en_reg_gen     : std_logic;
		    signal s_dut_uart_tx_i_data                : std_logic_vector(c_dut_data_length-1 downto 0);
		    signal s_dut_uart_tx_o_ready               : std_logic;
		    signal s_dut_uart_tx_o_done                : std_logic;
		    signal s_dut_uart_tx_o_line                : std_logic;
			signal s_dut_uart_tx_o_error               : std_logic_vector(7 downto 0);

		    -- =====================================================================================================================================================================
			-- 03.05.02.04. core_uart_rx
			-- =====================================================================================================================================================================			
		    signal s_dut_uart_rx_o_data_en : std_logic;
		    signal s_dut_uart_rx_o_data    : std_logic_vector(c_dut_data_length-1 downto 0);
		    signal s_dut_uart_rx_o_ready   : std_logic;
		    signal s_dut_uart_rx_o_done    : std_logic;
			signal s_dut_uart_rx_o_done_r  : std_logic;
			signal s_dut_uart_rx_o_done_re : std_logic;
		    signal s_dut_uart_rx_i_line    : std_logic;
			signal s_dut_uart_rx_o_error   : std_logic_vector(7 downto 0);

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.03. HOST
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.05.03.01. clock
			-- =====================================================================================================================================================================
            signal s_hst_i_clk : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.03.02. reset
			-- =====================================================================================================================================================================
	        signal s_hst_i_rst : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.03.03. core_uart_tx
			-- =====================================================================================================================================================================			
		    signal s_hst_uart_tx_i_data_en : std_logic;
		    signal s_hst_uart_tx_i_data_en_reg : std_logic_vector(c_ratio_clk_sim_clk_hst-1 downto 0);
			signal s_hst_uart_tx_i_data_en_reg_gen_tmp : std_logic_vector(c_ratio_clk_sim_clk_hst-1 downto 0);
			signal s_hst_uart_tx_i_data_en_reg_gen : std_logic;
		    signal s_hst_uart_tx_i_data    : std_logic_vector(c_hst_data_length-1 downto 0);
		    signal s_hst_uart_tx_o_ready   : std_logic;
		    signal s_hst_uart_tx_o_done    : std_logic;
		    signal s_hst_uart_tx_o_line    : std_logic;
			signal s_hst_uart_tx_o_error   : std_logic_vector(7 downto 0);

		    -- =====================================================================================================================================================================
			-- 03.05.03.04. core_uart_rx
			-- =====================================================================================================================================================================			
		    signal s_hst_uart_rx_o_data_en : std_logic;
		    signal s_hst_uart_rx_o_data    : std_logic_vector(c_hst_data_length-1 downto 0);
		    signal s_hst_uart_rx_o_ready   : std_logic;
		    signal s_hst_uart_rx_o_done    : std_logic;
			signal s_hst_uart_rx_o_done_r  : std_logic;
			signal s_hst_uart_rx_o_done_re : std_logic;
		    signal s_hst_uart_rx_i_line    : std_logic;
			signal s_hst_uart_rx_o_error   : std_logic_vector(7 downto 0);

begin

    -- =============================================================================================================================================================================
	-- 03.06. reset management
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_sim_rst <= '1','0' after c_sim_rst_delay;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. DUT
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_dut_i_rst <= '1','0' after c_dut_rst_delay;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.03. HOST
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_hst_i_rst <= '1','0' after c_hst_rst_delay;

    -- =============================================================================================================================================================================
	-- 03.07. clock generation
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_sim_clk : process
		begin
	        s_sim_clk <= '0';
	        wait for c_sim_clk_delay;
		    while true loop
		        s_sim_clk <= '1';
			    wait for c_sim_clk_period_ns/2;
			    s_sim_clk <= '0';
			    wait for c_sim_clk_period_ns/2;
		    end loop;
	    end process p_gen_sim_clk;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.02. oscillator
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_osc : process
		begin
	        s_osc <= '0';
	        wait for c_osc_delay;
		    while true loop
		        s_osc <= '1';
			    wait for c_osc_period_ns/2;
			    s_osc <= '0';
			    wait for c_osc_period_ns/2;
		    end loop;
	    end process p_gen_osc;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.03. HOST
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_hst_clk : process
		begin
	        s_hst_clk <= '0';
	        wait for c_hst_clk_delay;
		    while true loop
		        s_hst_clk <= '1';
			    wait for c_hst_clk_period_ns/2;
			    s_hst_clk <= '0';
			    wait for c_hst_clk_period_ns/2;
		    end loop;
	    end process p_gen_hst_clk;

    -- =============================================================================================================================================================================
	-- 03.08. clock assignment
    -- =============================================================================================================================================================================
    s_dut_i_clk <= s_osc;
	s_hst_i_clk <= s_hst_clk;

    -- =============================================================================================================================================================================
	-- 03.09. component instantiation
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.09.01. HOST : core_uart
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_hst_core_uart : core_uart
            generic map (
	             g_clk_i_freq  => c_hst_clk_freq
		        ,g_baud        => c_hst_baud
		        ,g_data_length => c_hst_data_length
	        )
            port map (
	             i_clk        => s_hst_i_clk
		        ,i_rst        => s_hst_i_rst
		        ,i_tx_data_en => s_hst_uart_tx_i_data_en_reg_gen
		        ,i_tx_data    => s_hst_uart_tx_i_data
		        ,o_tx_ready   => s_hst_uart_tx_o_ready
		        ,o_tx_done    => s_hst_uart_tx_o_done
		        ,o_tx_line    => s_hst_uart_tx_o_line
		        ,o_tx_error   => s_hst_uart_tx_o_error
		        ,o_rx_data_en => s_hst_uart_rx_o_data_en
		        ,o_rx_data    => s_hst_uart_rx_o_data
		        ,o_rx_ready   => s_hst_uart_rx_o_ready
		        ,o_rx_done    => s_hst_uart_rx_o_done
		        ,i_rx_line    => s_hst_uart_rx_i_line
		        ,o_rx_error   => s_hst_uart_rx_o_error
	        );

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.09.02. loopback
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_dut_uart_rx_i_line <= transport s_hst_uart_tx_o_line after 10 us;
		s_hst_uart_rx_i_line <= transport s_dut_uart_tx_o_line after 10 us;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.09.03. DUT : core_uart
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_dut_core_uart : core_uart
            generic map (
	             g_clk_i_freq  => c_dut_clk_freq
		        ,g_baud        => c_dut_baud
		        ,g_data_length => c_dut_data_length
	        )
            port map (
	             i_clk        => s_dut_i_clk
		        ,i_rst        => s_dut_i_rst
		        ,i_tx_data_en => s_dut_uart_tx_i_data_en_reg_gen
		        ,i_tx_data    => s_dut_uart_tx_i_data
		        ,o_tx_ready   => s_dut_uart_tx_o_ready
		        ,o_tx_done    => s_dut_uart_tx_o_done
		        ,o_tx_line    => s_dut_uart_tx_o_line
		        ,o_tx_error   => s_dut_uart_tx_o_error
		        ,o_rx_data_en => s_dut_uart_rx_o_data_en
		        ,o_rx_data    => s_dut_uart_rx_o_data
		        ,o_rx_ready   => s_dut_uart_rx_o_ready
		        ,o_rx_done    => s_dut_uart_rx_o_done
		        ,i_rx_line    => s_dut_uart_rx_i_line
		        ,o_rx_error   => s_dut_uart_rx_o_error
	        );

    -- =============================================================================================================================================================================
	-- 03.10. clock domain crossing (CDC)
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.10.01. from SIM to DUT (from fast to slow)
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_dut_uart_tx_i_data_en_sr: process(s_sim_rst,s_sim_clk)
		begin
		    if (s_sim_rst = '1') then
			    s_dut_uart_tx_i_data_en_reg <= (others => '0');
			elsif (rising_edge(s_sim_clk)) then
			    s_dut_uart_tx_i_data_en_reg <= s_dut_uart_tx_i_data_en_reg(s_dut_uart_tx_i_data_en_reg'length-2 downto 0) & s_dut_uart_tx_i_data_en;
			end if;
		end process s_dut_uart_tx_i_data_en_sr;
 
        s_dut_uart_tx_i_data_en_reg_gen_tmp(0) <= s_dut_uart_tx_i_data_en_reg(0);
		
		or_gen_dut_uart_tx_o_data_en : for i in 1 to c_ratio_clk_sim_clk_dut-1 generate
		    s_dut_uart_tx_i_data_en_reg_gen_tmp(i) <= s_dut_uart_tx_i_data_en_reg(i) or s_dut_uart_tx_i_data_en_reg_gen_tmp(i-1);
		end generate or_gen_dut_uart_tx_o_data_en;
		
		s_dut_uart_tx_i_data_en_reg_gen <= s_dut_uart_tx_i_data_en_reg_gen_tmp(s_dut_uart_tx_i_data_en_reg_gen_tmp'length-1);

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.10.02. from SIM to HST (from fast to slow)
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_hst_uart_tx_i_data_en_sr: process(s_sim_rst,s_sim_clk)
		begin
		    if (s_sim_rst = '1') then
			    s_hst_uart_tx_i_data_en_reg <= (others => '0');
			elsif (rising_edge(s_sim_clk)) then
			    s_hst_uart_tx_i_data_en_reg <= s_hst_uart_tx_i_data_en_reg(s_hst_uart_tx_i_data_en_reg'length-2 downto 0) & s_hst_uart_tx_i_data_en;
			end if;
		end process s_hst_uart_tx_i_data_en_sr;
 
        s_hst_uart_tx_i_data_en_reg_gen_tmp(0) <= s_hst_uart_tx_i_data_en_reg(0);
		
		or_gen_hst_uart_tx_o_data_en : for i in 1 to c_ratio_clk_sim_clk_hst-1 generate
		    s_hst_uart_tx_i_data_en_reg_gen_tmp(i) <= s_hst_uart_tx_i_data_en_reg(i) or s_hst_uart_tx_i_data_en_reg_gen_tmp(i-1);
		end generate or_gen_hst_uart_tx_o_data_en;
		
		s_hst_uart_tx_i_data_en_reg_gen <= s_hst_uart_tx_i_data_en_reg_gen_tmp(s_hst_uart_tx_i_data_en_reg_gen_tmp'length-1);
			
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.10.03. edge detector from HST to SIM (from slow to fast) 
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		p_hst_uart_rx_o_done_re : process(s_sim_rst,s_sim_clk)
        begin
		    if (s_sim_rst = '1') then
			    s_hst_uart_rx_o_done_r <= '0';
				s_hst_uart_rx_o_done_re <= '0';
			elsif (rising_edge(s_sim_clk)) then
			    s_hst_uart_rx_o_done_r <= s_hst_uart_rx_o_done;
				if (s_hst_uart_rx_o_done = '1' and s_hst_uart_rx_o_done_r = '0') then
				    s_hst_uart_rx_o_done_re <= '1';
				else
				    s_hst_uart_rx_o_done_re <= '0';
				end if;
			end if;
        end process p_hst_uart_rx_o_done_re;	
			
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.10.04. edge detector from DUT to SIM (from slow to fast) 
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		p_dut_uart_rx_o_done_re : process(s_sim_rst,s_sim_clk)
        begin
		    if (s_sim_rst = '1') then
			    s_dut_uart_rx_o_done_r <= '0';
				s_dut_uart_rx_o_done_re <= '0';
			elsif (rising_edge(s_sim_clk)) then
			    s_dut_uart_rx_o_done_r <= s_dut_uart_rx_o_done;
				if (s_dut_uart_rx_o_done = '1' and s_dut_uart_rx_o_done_r = '0') then
				    s_dut_uart_rx_o_done_re <= '1';
				else
				    s_dut_uart_rx_o_done_re <= '0';
				end if;
			end if;
        end process p_dut_uart_rx_o_done_re;
			
    -- =============================================================================================================================================================================
	-- 03.11. fsm_main
    -- =============================================================================================================================================================================
	p_fsm_main : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_main_state <= state_fsm_main_start;
			s_sim_done <= '0';
			s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_done <= '0';
            s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
		    case s_fsm_main_state is
			    -- wait for DUT reset deassertion
				when state_fsm_main_start =>
				    if (s_dut_i_rst = '0') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_open;
						s_sim_file_req_rpt_open <= '1';
					end if;
				-- wait for RPT file to be opened
			    when state_fsm_main_file_rpt_open =>
				    if (s_sim_file_ack_rpt_open = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_open;
					    s_sim_file_req_log_open <= '1';
					end if;
				-- wait for LOG file to be opened
				when state_fsm_main_file_log_open =>
				    if (s_sim_file_ack_log_open = '1') then
					    s_fsm_main_state <= state_fsm_main_init;
						s_sim_init_req <= '1';
					end if;
				-- waiting for init done
				when state_fsm_main_init =>
				    if (s_sim_init_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_run;
						-- run test
					    s_sim_test_req <= '1';
					end if;
				-- waiting for test done
				when state_fsm_main_run =>
                    if (s_sim_test_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_close;
						s_sim_file_req_log_close <= '1';
					end if;
				-- waiting for data file to be closed
				when state_fsm_main_file_log_close =>
                    if (s_sim_file_ack_log_close = '1') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_close;
						s_sim_file_req_rpt_close <= '1';
					end if;
				-- waiting for SIM report file to be closed
				when state_fsm_main_file_rpt_close =>
                    if (s_sim_file_ack_rpt_close = '1') then
					    s_fsm_main_state <= state_fsm_main_stop;
				        s_sim_done <= '1';
					end if;
				-- test stopped
                when state_fsm_main_stop =>
                    null;
			end case;
		end if;
	end process p_fsm_main;

    -- =============================================================================================================================================================================
	-- 03.12. fsm_init
    -- =============================================================================================================================================================================
	fsm_init : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_init_state <= state_fsm_init_idle;
			s_sim_init_ack <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_init_ack <= '0';
		    case s_fsm_init_state is
			    -- waiting for init request
			    when state_fsm_init_idle =>
				    if (s_sim_init_req = '1') then
					    s_fsm_init_state <= state_fsm_init_run;
					end if;
				-- running init
				when state_fsm_init_run =>
					s_fsm_init_state <= state_fsm_init_done;
                    s_sim_init_ack <= '1';
				-- init done
                when state_fsm_init_done =>
				    null;
			end case;
		end if;
	end process fsm_init;

    -- =============================================================================================================================================================================
	-- 03.13. fsm_test
    -- =============================================================================================================================================================================
	p_fsm_test : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
			s_sim_test_ack <= '0';
			s_dut_uart_tx_i_data_en <= '0';
			s_dut_uart_tx_i_data <= (others => '0');
			s_hst_uart_tx_i_data_en <= '0';
			s_hst_uart_tx_i_data <= (others => '0');
			s_array_data_cnt <= 0;
			s_sim_test_status <= TEST_OK;
			s_error_test <= '0';
		    s_fsm_test_state <= state_fsm_test_idle;
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_test_ack <= '0';
		    case s_fsm_test_state is
			    -- waiting for test request
			    when state_fsm_test_idle =>
				    if (s_sim_test_req = '1') then
					    s_fsm_test_state <= state_fsm_test_dut_to_hst_send_data;
					end if;
                -- send data to HOST uart receiver
                when state_fsm_test_dut_to_hst_send_data =>
                    s_dut_uart_tx_i_data <= c_array_data(s_array_data_cnt);
                    s_dut_uart_tx_i_data_en <= '1';
					s_fsm_test_state <= state_fsm_test_dut_to_hst_wait_ready;
				when state_fsm_test_dut_to_hst_wait_ready =>
                    s_dut_uart_tx_i_data_en <= '0';
					s_fsm_test_state <= state_fsm_test_dut_to_hst_wait_done;
                when state_fsm_test_dut_to_hst_wait_done =>
				    -- data received
				    if (s_hst_uart_rx_o_done_re = '1') then
					    s_fsm_test_state <= state_fsm_test_dut_to_hst_check_data;
					end if;
                when state_fsm_test_dut_to_hst_check_data =>
				    if (s_hst_uart_rx_o_data_en = '1') then
					    -- error detection
					    if (s_hst_uart_rx_o_data /= c_array_data(s_array_data_cnt)) then
						    s_error_test <= '1';
							s_array_data_cnt <= 0;
							s_sim_test_ack <= '1';
							s_sim_test_status <= TEST_KO;
							s_fsm_test_state <= state_fsm_test_done;
						-- data received is valid
                        else
						    -- all data transmitted
						    if (s_array_data_cnt = c_array_data_length-1) then
							    s_array_data_cnt <= 0;
								s_fsm_test_state <= state_fsm_test_hst_to_dut_send_data;
							else
						        s_array_data_cnt <= s_array_data_cnt + 1;
							    s_fsm_test_state <= state_fsm_test_dut_to_hst_send_data;

							end if;
						end if;
					end if;
                -- send data to DUT uart receiver
                when state_fsm_test_hst_to_dut_send_data =>
                    s_hst_uart_tx_i_data <= c_array_data(s_array_data_cnt);
                    s_hst_uart_tx_i_data_en <= '1';
					s_fsm_test_state <= state_fsm_test_hst_to_dut_wait_ready;
				when state_fsm_test_hst_to_dut_wait_ready =>
                    s_hst_uart_tx_i_data_en <= '0';
                    s_fsm_test_state <= state_fsm_test_hst_to_dut_wait_done;
                when state_fsm_test_hst_to_dut_wait_done =>
				    -- data received
				    if (s_dut_uart_rx_o_done_re = '1') then
					    s_fsm_test_state <= state_fsm_test_hst_to_dut_check_data;
					end if;
                when state_fsm_test_hst_to_dut_check_data =>
				    if (s_dut_uart_rx_o_data_en = '1') then
					    -- error detection
					    if (s_dut_uart_rx_o_data /= c_array_data(s_array_data_cnt)) then
						    s_error_test <= '1';
							s_array_data_cnt <= 0;
							s_sim_test_ack <= '1';
							s_sim_test_status <= TEST_KO;
							s_fsm_test_state <= state_fsm_test_done;
						-- data received is valid
                        else
						    -- all data transmitted
						    if (s_array_data_cnt = c_array_data_length-1) then
							    s_array_data_cnt <= 0;
							    s_sim_test_ack <= '1';
							    s_sim_test_status <= TEST_OK;
								s_fsm_test_state <= state_fsm_test_done;
							else
						        s_array_data_cnt <= s_array_data_cnt + 1;
							    s_fsm_test_state <= state_fsm_test_hst_to_dut_send_data;
							end if;
						end if;
					end if;
				-- test done
                when state_fsm_test_done =>
                    null;
			end case;
		end if;
	end process p_fsm_test;

    -- =============================================================================================================================================================================
	-- 03.14. fsm_file_mgt_log
    -- =============================================================================================================================================================================
	p_fsm_file_mgt_log : process(s_sim_rst,s_sim_clk)
		constant c_justified  : side   := right;
		constant c_field      : width  := 0;
		constant c_unit       : time   := ns;
		constant c_separator  : string := ",";
		constant c_value_head : string := "time,data";
	    variable v_value_time : time;
		variable v_value_data : string(1 to 4);
		variable v_value_foot : string(1 to 7);
		variable v_line       : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_open;
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
            case s_fsm_file_mgt_log is
                -- open file
			    when state_fsm_file_mgt_log_open =>
				    if (s_sim_file_req_log_open = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_head;
						s_sim_file_ack_log_open <= '1';
						proc_file_log_open(c_file_log_name,f_file_log);
					end if;
				-- write header
				when state_fsm_file_mgt_log_write_head =>
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_data;
						write(v_line,c_value_head,c_justified,c_field);
	                    writeline(f_file_log,v_line);
				-- write data
				when state_fsm_file_mgt_log_write_data =>
				    if (s_sim_file_req_log_close = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_close;
						-- timestamp
						v_value_time := now;
						write(v_line,v_value_time,c_justified,c_field,c_unit);
						-- separator
						write(v_line,c_separator,c_justified,c_field);
						-- data value
						v_value_data := "NONE";
					    write(v_line,v_value_data,c_justified,c_field);
	                    writeline(f_file_log,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_log_close =>
					s_fsm_file_mgt_log <= state_fsm_file_mgt_log_done;
				    s_sim_file_ack_log_close <= '1';
                    proc_file_log_close(c_file_log_name,f_file_log);
				-- done
				when state_fsm_file_mgt_log_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_log;

    -- =============================================================================================================================================================================
	-- 03.15. fsm_file_mgt_rpt
    -- =============================================================================================================================================================================
	p_fsm_file_mgt_rpt : process(s_sim_rst,s_sim_clk)
		constant c_justified    : side  := right;
		constant c_field        : width := 0;
		variable v_value_status : string(1 to 7);
		variable v_line         : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_open;
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
            case s_fsm_file_mgt_rpt is
                -- open file
			    when state_fsm_file_mgt_rpt_open =>
				    if (s_sim_file_req_rpt_open = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_write_status;
						s_sim_file_ack_rpt_open <= '1';
						proc_file_rpt_open(c_file_rpt_name,f_file_rpt);
					end if;
				-- write status
				when state_fsm_file_mgt_rpt_write_status =>
				    if (s_sim_file_req_rpt_close = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_close;
					    -- write test status
					    case s_sim_test_status is
					        when TEST_OK => v_value_status := "TEST_OK";
						    when others  => v_value_status := "TEST_KO";
					    end case;
					    write(v_line,v_value_status,c_justified,c_field);
	                    writeline(f_file_rpt,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_rpt_close =>
					s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_done;
				    s_sim_file_ack_rpt_close <= '1';
                    proc_file_rpt_close(c_file_rpt_name,f_file_rpt);
				-- done
				when state_fsm_file_mgt_rpt_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_rpt;

    -- =============================================================================================================================================================================
	-- 03.16. error detection
    -- =============================================================================================================================================================================
	p_check_dut_error : process(s_dut_i_rst,s_sim_clk)
	    variable v_error : std_logic;
	begin
	    if (s_dut_i_rst = '1') then
	        v_error := '0';
			s_error <= '0';
	    elsif (rising_edge(s_sim_clk)) then
		    v_error := '0';
			-- parsing error vector
		    for i in 0 to s_dut_uart_tx_o_error'length-1 loop
		        -- error detected
			    if (s_dut_uart_tx_o_error(i) = '1') then
				    v_error := '1';
				end if;
			end loop;
			s_error <= v_error;
		end if;
	end process p_check_dut_error;	
	
    -- =============================================================================================================================================================================
	-- 03.17. simulation abort
    -- =============================================================================================================================================================================
	p_sim_abort : process(s_sim_clk)
	begin
		if (rising_edge(s_sim_clk)) then
            if (s_error = '1') then
			    assert false 
				    report "end of simulation - DUT error detected" 
					    severity failure;
			end if;
			if (s_error_test = '1') then
			    assert false 
				    report "end of simulation - Test error detected" 
					    severity failure;
			end if;
		end if;
	end process p_sim_abort;

    -- =============================================================================================================================================================================
	-- 03.18. end of simulation
    -- =============================================================================================================================================================================
	p_sim_end : process(s_sim_clk)
	begin
		if (rising_edge(s_sim_clk)) then
            if (s_sim_done = '1') then
			    assert false 
				    report "end of simulation - success" 
					    severity failure;
			end if;
		end if;
	end process p_sim_end;

end architecture behavioral;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################