-- #################################################################################################################################################################################
-- file :
--     core_uart_tx.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     UART transmitter
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     register tranfer level (RTL)
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     clock ratio must be higher or equal to 16.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2024-04-23
--         file creation
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--     02. entity
--     03. architecture
--         03.01. constants
--         03.02. signals
--         03.03. input assignment
--         03.04. alive output pin generation
--         03.05. output assignment
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;

    -- =============================================================================================================================================================================
	-- 01.01. custom
    -- =============================================================================================================================================================================	
	library work;
	    use work.pkg_core_uart_tx.all;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity core_uart_tx is
    generic (
	     g_clk_i_freq  : integer := 100_000_000
		;g_baud        : integer :=     115_200
		;g_data_length : integer :=           8
	);
    port (
	     i_clk     : in  std_logic
		;i_rst     : in  std_logic
		;i_data_en : in  std_logic
		;i_data    : in  std_logic_vector(g_data_length-1 downto 0)
		;o_ready   : out std_logic
		;o_done    : out std_logic
		;o_tx      : out std_logic
		;o_error   : out std_logic_vector(7 downto 0)
	);
end entity core_uart_tx;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture rtl of core_uart_tx is

    -- =============================================================================================================================================================================
	-- 03.01. constants
    -- =============================================================================================================================================================================
	constant c_clk_ratio : integer := integer(real(g_clk_i_freq)/real(g_baud));

    -- =============================================================================================================================================================================
	-- 03.04. types
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. FSM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        type t_fsm_main is (
		     state_fsm_main_idle
		    ,state_fsm_main_start
			,state_fsm_main_data
			,state_fsm_main_stop
		);
	
    -- =============================================================================================================================================================================
	-- 03.02. signals
    -- =============================================================================================================================================================================
	signal s_clk         : std_logic;
	signal s_rst         : std_logic;
	signal s_error_ratio : std_logic;
	signal s_data        : std_logic_vector(g_data_length-1 downto 0);
	signal s_data_en     : std_logic;
	signal s_data_reg    : std_logic_vector(g_data_length-1 downto 0);
	signal s_cnt_clk     : integer range 0 to c_clk_ratio-1;
	signal s_cnt_bit     : integer range 0 to g_data_length-1;
	signal s_tx          : std_logic;
	signal s_ready       : std_logic;
	signal s_done        : std_logic;
	signal s_fsm_main    : t_fsm_main;
	
begin
    -- =============================================================================================================================================================================
	-- 03.03. check input parameters
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. check clock ratio
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    check_clk_ratio_ok : if (c_clk_ratio > c_clk_ratio_upper_bound or c_clk_ratio = c_clk_ratio_upper_bound) generate
	        s_error_ratio <= '0';
	    end generate check_clk_ratio_ok;

	    check_clk_ratio_ko : if (c_clk_ratio < c_clk_ratio_upper_bound) generate
	        s_error_ratio <= '1';
	    end generate check_clk_ratio_ko;

    -- =============================================================================================================================================================================
	-- 03.04. input assignment
    -- =============================================================================================================================================================================
	s_clk     <= i_clk;
	s_rst     <= i_rst;
    s_data    <= i_data;
	s_data_en <= i_data_en;

    -- =============================================================================================================================================================================
	-- 03.05. main FSM
    -- =============================================================================================================================================================================
    p_fsm_main : process(s_clk,s_rst)
	begin
	    if (s_rst = '1') then
		    s_data_reg <= (others => '0');
			s_cnt_clk <= 0;
			s_cnt_bit <= 0;
			s_tx <= '1';
			s_ready <= '1';
			s_done  <= '0';
			s_fsm_main <= state_fsm_main_idle;
		elsif (rising_edge(s_clk)) then
		    s_done <= '0';
		    case s_fsm_main is
			    when state_fsm_main_idle =>
				    s_ready <= '1';
				    if (s_data_en = '1') then
					    s_ready <= '0';
					    s_data_reg <= s_data;
					    s_fsm_main <= state_fsm_main_start;
					end if;
				when state_fsm_main_start =>
				    -- start bit
				    s_tx <= '0';
				    if (s_cnt_clk = c_clk_ratio-1) then
					    s_cnt_clk <= 0;
						s_fsm_main <= state_fsm_main_data;
					else
					    s_cnt_clk <= s_cnt_clk + 1;
					end if;
				when state_fsm_main_data  =>
				    s_tx <= s_data_reg(s_data_reg'high);
				    if (s_cnt_clk = c_clk_ratio-1) then
					    s_cnt_clk <= 0;
						-- shifting data to the right
						s_data_reg <= s_data_reg(g_data_length-2 downto 0) & '0';
						if (s_cnt_bit =  g_data_length-1) then
						    s_cnt_bit <= 0;
						    s_fsm_main <= state_fsm_main_stop;
						else
						    -- transmitting next data bit
						    s_cnt_bit <= s_cnt_bit + 1;
						end if;
					else
					    s_cnt_clk <= s_cnt_clk + 1;
					end if;
				when state_fsm_main_stop  =>
				    -- stop bit
				    s_tx <= '1';
				    if (s_cnt_clk = c_clk_ratio-1) then
					    s_cnt_clk <= 0;
						s_ready <= '1';
						s_done <= '1';
						s_fsm_main <= state_fsm_main_idle;
					else
					    s_cnt_clk <= s_cnt_clk + 1;
					end if;
			end case;
		end if;
	end process p_fsm_main;

    -- =============================================================================================================================================================================
	-- 03.06. output assignment
    -- =============================================================================================================================================================================
	o_done  <= s_done;
	o_tx    <= s_tx;
	o_ready <= s_ready;
    o_error <= (
	     c_pos_error_ratio => s_error_ratio
		,others            => '0'
	);

end architecture rtl;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################